module ALU_tb;
  reg [31:0] a,b;
  reg [2:0] opcode;
  wire [63:0] res;
  wire ov;
  
  ALU DUT(.a(a), .b(b), .opcode(opcode), .res(res), .ov(ov));
  
  initial
    begin
      a = 32'b00000000000000000000000000000001;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b000;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000101;
      opcode = 3'b001;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b010;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b011;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b100;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b101;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b110;
      #10;
      
      a = 32'b00000000000000000000000000001111;
      b = 32'b00000000000000000000000000000010;
      opcode = 3'b111;
      #10;
      
      $finish;
    end
endmodule